module fifo(
	// write interface
	clk_i, rst_i, wdata_i, wr_en_i, wr_error_o,
	// read interface	
	rdata_o, full_o, empty_o, rd_en_i, rd_error_o
	
);

parameter DEPTH=16, WIDTH=8, PTR_WIDTH=4;

//wr_ptr is internal to the design 
input clk_i, rst_i, wr_en_i, rd_en_i;
input [WIDTH-1:0] wdata_i;
output reg wr_error_o, rd_error_o, full_o, empty_o;
output reg [WIDTH-1:0] rdata_o;

// mem declaration 
reg [WIDTH-1:0] mem [DEPTH-1:0];

// internal signals
reg [PTR_WIDTH-1:0] rd_ptr, wr_ptr;
reg wr_toggle_f, rd_toggle_f;

integer i; // Remember to remove unwanted integers

always @(posedge clk_i) begin 
	if (rst_i == 1) begin 
		wr_error_o = 0;
		rd_error_o = 0;
		full_o = 0;
		empty_o = 1;
		rdata_o = 0;
		rd_ptr = 0;
		wr_ptr = 0;
		wr_toggle_f = 0;
		rd_toggle_f = 0;
		// clear the memory
		for (i=0; i<DEPTH; i=i+1) begin 
			mem[i] = 0;	
		end
	end	

	else begin 
		wr_error_o = 0;
		rd_error_o = 0;
		if (wr_en_i == 1) begin 
			if (full_o == 1) begin 
				wr_error_o = 1;
			end 
			else begin 
				// store data into memory
				mem[wr_ptr] = wdata_i;
				// increment the wr_ptr
				if (wr_ptr == DEPTH-1) wr_toggle_f = ~wr_toggle_f;
				wr_ptr = wr_ptr + 1;
			end
		end

		if (rd_en_i == 1) begin
			if (empty_o == 1) begin 
				rd_error_o = 1;
			end
			else begin 
				rdata_o = mem[rd_ptr];
				// increment the rd_ptr
				if (rd_ptr == DEPTH-1) rd_toggle_f = ~rd_toggle_f;
				rd_ptr = rd_ptr + 1;
			end 		
		end
	end 
end 



// logic to create empty and full condition

always @(*) begin 
	empty_o = 0;
	full_o = 0;
	if (rd_ptr == wr_ptr) begin 
		if (wr_toggle_f == rd_toggle_f) empty_o = 1;
		if (wr_toggle_f != rd_toggle_f) full_o = 1;		
	end
end

endmodule


